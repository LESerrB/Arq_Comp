library verilog;
use verilog.vl_types.all;
entity logint_vlg_vec_tst is
end logint_vlg_vec_tst;
