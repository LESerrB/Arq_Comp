library verilog;
use verilog.vl_types.all;
entity reg_mpc_vlg_vec_tst is
end reg_mpc_vlg_vec_tst;
