library verilog;
use verilog.vl_types.all;
entity increm_vlg_vec_tst is
end increm_vlg_vec_tst;
