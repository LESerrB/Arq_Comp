library verilog;
use verilog.vl_types.all;
entity mem_vlg_vec_tst is
end mem_vlg_vec_tst;
