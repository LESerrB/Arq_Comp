library verilog;
use verilog.vl_types.all;
entity interr_trans_vlg_vec_tst is
end interr_trans_vlg_vec_tst;
