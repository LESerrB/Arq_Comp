library verilog;
use verilog.vl_types.all;
entity muxdir_vlg_vec_tst is
end muxdir_vlg_vec_tst;
