library verilog;
use verilog.vl_types.all;
entity logsel_vlg_check_tst is
    port(
        CC              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end logsel_vlg_check_tst;
