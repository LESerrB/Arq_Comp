library verilog;
use verilog.vl_types.all;
entity secuen_completo_vlg_vec_tst is
end secuen_completo_vlg_vec_tst;
