library verilog;
use verilog.vl_types.all;
entity logsel_vlg_vec_tst is
end logsel_vlg_vec_tst;
