library verilog;
use verilog.vl_types.all;
entity registrosmemoria_vlg_vec_tst is
end registrosmemoria_vlg_vec_tst;
